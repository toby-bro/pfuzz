module buf_primitive (
    input wire i,
    output wire o
);
    buf b1 (o, i);
endmodule

