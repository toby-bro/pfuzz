module mod_default_disable (
    input bit enable_in,
    output bit out
);
    assign out = enable_in;
endmodule

