module ConcatVectorOps (
    input logic [3:0] a,
    input logic [3:0] b,
    input logic [7:0] c,
    output logic [15:0] out_concat
);
    assign out_concat = {a, b, c};
endmodule

