module generic_class_scope_diag_mod (
    input logic [7:0] in_val,
    output logic [7:0] out_val
);
    assign out_val = in_val;
endmodule

