module bind_module (
    input logic bind_in,
    output logic bind_out
);
    assign bind_out = bind_in;
endmodule

