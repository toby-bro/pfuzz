module another_module_config_dummy (
    input logic i,
    output logic o
);
 assign o = i & i; 
endmodule

