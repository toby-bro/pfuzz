module configuration_top (
    input logic i_in,
    output logic o_out
);
    assign o_out = i_in;
endmodule

