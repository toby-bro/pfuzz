module DummyHierModule (
    input bit in_bit,
    output logic out_logic
);
    assign out_logic = in_bit;
endmodule

