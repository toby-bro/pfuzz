module ImplicitTimeScaleModule (
    input logic in_its,
    output logic out_its
);
    assign out_its = in_its;
endmodule

