module WiredNet (
	data1,
	data2,
	out_wired
);
	input wire data1;
	input wire data2;
	output wire out_wired;
	wor w_or;
	assign w_or = data1;
	assign w_or = data2;
	assign out_wired = w_or;
endmodule