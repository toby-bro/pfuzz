module child_empty_ports (
    p1,
    p2
);
    input logic p1;
    output logic p2;
    assign p2 = p1;
endmodule

