module ModuleBasicDisplay(
    input wire [7:0] data_in,
    input wire enable,
    output reg [7:0] data_out
);
always @* begin
    data_out = data_in;
    if (enable) begin
        $display("ModuleBasicDisplay: data_in = %d", data_in);
        $write("ModuleBasicDisplay: data_in = %h\n", data_in);
        $displayb("Binary data_in: %b", data_in);
        $displayo("Octal data_in: %o", data_in);
        $displayh("Hex data_in: %h", data_in);
        $writeb("Binary data_in: %b\n", data_in);
        $writeo("Octal data_in: %o\n", data_in);
        $writeh("Hex data_in: %h\n", data_in);
        $display("Multiple args: %d %h %b", data_in, data_in, data_in);
    end
end
endmodule
module ModuleMonitorStrobe(
    input wire [7:0] data_in_monitor,
    input wire clk_monitor,
    input wire enable_monitor,
    output reg [7:0] data_out_monitor
);
always @(posedge clk_monitor) begin
    data_out_monitor <= data_in_monitor;
    if (enable_monitor) begin
        $monitor("ModuleMonitorStrobe: data_in=%d data_out=%d", data_in_monitor, data_out_monitor);
        $monitorb("Monitor Binary: %b", data_in_monitor);
        $monitoro("Monitor Octal: %o", data_in_monitor);
        $monitorh("Monitor Hex: %h", data_in_monitor);
    end
end
always @* begin
    if (enable_monitor && data_in_monitor > 100) begin
       $strobe("ModuleMonitorStrobe: Strobe! data_in=%d data_out=%d", data_in_monitor, data_out_monitor);
       $strobeb("Strobe Binary: %b", data_in_monitor);
       $strobeo("Strobe Octal: %o", data_in_monitor);
       $strobeh("Strobe Hex: %h", data_in_monitor);
    end
end
endmodule
module ModuleSeverity(
    input wire [3:0] level_severity,
    input wire enable_severity,
    output reg dummy_out_severity
);
always @* begin
    dummy_out_severity = enable_severity;
    if (enable_severity) begin
        $info("ModuleSeverity: Info message with data %0d", level_severity);
        $warning("ModuleSeverity: Warning message with data %0d", level_severity);
        $error("ModuleSeverity: Error message with data %0d", level_severity);
        case (level_severity)
            0: $fatal(0);
            1: $fatal(1, "ModuleSeverity: Fatal message with code %0d and data %0d", 1, level_severity);
            default: ;
        endcase
    end
end
endmodule
module ModuleFileIO(
    input wire [7:0] data_in_file,
    input wire enable_file,
    output reg dummy_out_file
);
integer file_handle;
reg [7:0] memory [0:7];
reg [15:0] wide_memory [0:3];
string string_memory [0:3];
string sreadmem_str;
reg [31:0] sreadmem_dummy_output; 
always @* begin
    dummy_out_file = enable_file;
    file_handle = 32'h8000_0001; 
    if (enable_file) begin
        $fdisplay(file_handle, "ModuleFileIO: Data in file: %0d", data_in_file);
        $fwrite(file_handle, "ModuleFileIO: Data in file (hex): %h\n", data_in_file);
        $fdisplayb(file_handle, "File Binary: %b", data_in_file);
        $fwriteo(file_handle, "File Octal: %o\n", data_in_file);
        $fdisplayh(file_handle, "File Hex: %h", data_in_file);
        $fwriteb(file_handle, "File Binary: %b\n", data_in_file);
        $readmemb("dummy.mem", memory);
        $readmemh("dummy_wide.mem", wide_memory, 0, 3);
        $writememb("output.mem", memory);
        $writememh("output_wide.mem", wide_memory, 1, 2);
        string_memory[0] = "abc"; string_memory[1] = "def"; string_memory[2] = "ghi"; string_memory[3] = "jkl";
        memory[0] = 8'h11; memory[1] = 8'h22; memory[2] = 8'h33; memory[3] = 8'h44;
        wide_memory[0] = 16'h1122; wide_memory[1] = 16'h3344; wide_memory[2] = 16'h5566; wide_memory[3] = 16'h7788;
        sreadmem_str = string_memory[0];
        $sreadmemb(memory, 0, 3, string_memory[0]);
        $sreadmemh(wide_memory, 0, 1, sreadmem_str);
        $sreadmemb(memory, 0, 7, "0123456789abcdef"); 
        $sreadmemh(wide_memory, 0, 3, "0123456789abcdef"); 
        $sreadmemh(wide_memory, 0, 3, "01234567", "89abcdef"); 
    end
end
endmodule
module ModuleStringOps(
    input wire [7:0] data_in_string,
    input wire enable_string,
    output string output_string
);
string format_string;
always @* begin
    output_string = "";
    format_string = "";
    if (enable_string) begin
        $swrite(output_string, "Data in string: %0d", data_in_string);
        $swriteb(output_string, " Data bin: %b", data_in_string);
        $swriteo(output_string, " Data oct: %o", data_in_string);
        $swriteh(output_string, " Data hex: %h", data_in_string);
        $sformat(format_string, "Formatted data: %b", data_in_string);
        $sformat(format_string, "Formatted data: %s %h", "Value", data_in_string);
        output_string = {output_string, " ", format_string};
    end
end
endmodule
module ModuleSystemCast(
    input wire [15:0] data_in_sc,
    input wire enable_sc,
    output reg [7:0] data_out_sc,
    output reg cast_success_sc
);
integer system_ret_val;
reg [7:0] cast_target;
always @* begin
    data_out_sc = data_in_sc[7:0];
    cast_success_sc = 0;
    if (enable_sc) begin
        system_ret_val = $system("echo 'test $system'");
        cast_success_sc = $cast(cast_target, data_in_sc);
        data_out_sc = cast_target;
    end
end
endmodule
module ModuleHierarchyTasks( 
    input wire hierarchy_in,
    input wire clk_hierarchy,
    input wire enable_hierarchy,
    output wire hierarchy_out
);
    assign hierarchy_out = hierarchy_in;
    reg hierarchy_var = 1'b0;
    always @(hierarchy_in) begin
        hierarchy_var = hierarchy_in;
    end
    always @(posedge clk_hierarchy) begin
        if (enable_hierarchy) begin
            $printtimescale; 
            $dumpvars; 
            $dumpvars(1); 
            $dumpvars(1, hierarchy_var); 
            $dumpports; 
            $sdf_annotate("timing.sdf");
            $assertcontrol(1, 1, 1, 1); 
            $asserton; 
            $assertoff; 
            $assertkill; 
            $assertpasson; 
            $assertpassoff; 
            $assertfailon; 
            $assertfailoff; 
            $assertnonvacuouson; 
            $assertvacuousoff; 
        end
    end
endmodule
module ModuleStochastic(
    input wire [31:0] seed1,
    input wire [31:0] seed2,
    input wire [31:0] seed3,
    input wire [31:0] add_item_in,
    input wire [31:0] add_weight_in,
    input wire [31:0] exam_index_in,
    input wire enable_stochastic,
    output reg [31:0] q_handle_out,
    output reg [31:0] q_item_out,
    output reg [31:0] q_weight_out,
    output reg [31:0] q_status_out
);
integer q_handle;
integer add_success;
integer removed_item, removed_weight, removed_status;
integer exam_item, exam_weight;
integer is_full_var;
integer dummy_output_qfull; 
always @* begin
    q_handle_out = 0;
    q_item_out = 0;
    q_weight_out = 0;
    q_status_out = 0;
    if (enable_stochastic) begin
        $q_initialize(seed1, seed2, seed3, q_handle);
        q_handle_out = q_handle;
        $q_add(q_handle, add_item_in, add_weight_in, add_success);
        q_status_out = add_success; 
        $q_remove(q_handle, removed_item, removed_weight, removed_status);
        q_item_out = removed_item; 
        q_weight_out = removed_weight;
        $q_exam(q_handle, exam_index_in, exam_item, exam_weight);
        q_item_out = exam_item;
        q_weight_out = exam_weight;
        is_full_var = $q_full(q_handle, dummy_output_qfull);
        q_status_out = is_full_var; 
    end
end
endmodule
module ModuleSimpleTasks(
    input wire [31:0] int_arg1,
    input string string_arg1,
    input wire enable_simple,
    output reg dummy_out_simple
);
integer system_ret_val; 
integer reset_arg1 = 1, reset_arg2 = 0, reset_arg3 = 1; 
always @* begin
    dummy_out_simple = enable_simple;
    system_ret_val = 0; 
    if (enable_simple) begin
        $timeformat(-9, 1, "ns", 0);
        $monitoron;
        $monitoroff;
        $dumpfile("vcd.vcd");
        $dumpon;
        $dumpoff;
        $dumpall;
        $dumplimit(int_arg1);
        $dumpflush;
        $dumpportson("dumpports.vcd");
        $dumpportsoff("dumpports.vcd");
        $dumpportsall("dumpports.vcd");
        $dumpportslimit(int_arg1, "dumpports.vcd");
        $dumpportsflush("dumpports.vcd");
        $input(string_arg1);
        $key(string_arg1);
        $key;
        $nokey;
        $log(string_arg1);
        $nolog;
        $reset(reset_arg1, reset_arg2, reset_arg3);
        $save("checkpoint.save");
        $restart("checkpoint.save");
        $incsave("inc_checkpoint.save");
        $showscopes(int_arg1);
        system_ret_val = $system(string_arg1); 
    end
end
endmodule
module ModuleStaticAssert(
    input wire input_val,
    output reg dummy_out_sa
);
    parameter STATIC_COND_TRUE = 1;
    parameter STATIC_COND_FALSE = 0;
    $static_assert(STATIC_COND_TRUE);
    $static_assert(STATIC_COND_TRUE, "Static assertion passed (True)");
    $static_assert(STATIC_COND_TRUE, "Static assertion passed with value %0d", STATIC_COND_TRUE);
    always @* begin
        dummy_out_sa = input_val;
    end
endmodule
module ModuleFinishStop(
    input wire enable_fs,
    input wire [7:0] status_fs,
    output reg dummy_out_fs
);
    always @* begin
        dummy_out_fs = enable_fs;
        if (enable_fs) begin
            $finish;
            $finish(status_fs); 
            $stop;
            $stop(status_fs); 
        end
    end
endmodule
