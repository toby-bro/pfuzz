module super_outside_class_diag_mod (
    input int in_val,
    output int out_val
);
    assign out_val = in_val;
endmodule

