module BindSimpleModule (
    input bit in,
    output bit out
);
    assign out = in;
endmodule

