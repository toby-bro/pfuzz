module net_var_conn_child (
    input logic in_logic,
    output logic out_wire
);
    assign out_wire = in_logic;
endmodule

