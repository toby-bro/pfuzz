module ModuleDefinition (
    input wire in_md,
    output logic out_md
);
    assign out_md = in_md;
endmodule

