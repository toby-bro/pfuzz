module mod_large_array_target (
    input logic in_la,
    output logic out_la
);
    assign out_la = in_la;
endmodule

