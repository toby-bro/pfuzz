module cu_base (
    input logic [7:0] data_in,
    output logic [7:0] data_out
);
    assign data_out = data_in;
endmodule

