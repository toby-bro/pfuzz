module ProgramDefinition (
    input wire in_pd,
    output logic out_pd
);
    assign out_pd = in_pd;
endmodule

