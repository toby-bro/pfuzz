module child_module_v2_config_dummy (
    input logic i,
    output logic o
);
 assign o = i | i; 
endmodule

