module explicit_non_ansi_decl_module (
    p_in,
    p_out
);
    input logic p_in;
    output wire p_out;
    assign p_out = p_in;
endmodule

