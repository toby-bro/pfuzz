module mod_simple (
    input wire in,
    output wire out
);
    assign out = in;
endmodule

