module module_using_package_param (
    input logic [31:0] wide_data_in,
    output logic [31:0] wide_data_out
);
    assign wide_data_out = wide_data_in;
endmodule

