module child_module_v1_config_dummy (
    input logic i,
    output logic o
);
 assign o = ~i; 
endmodule

