module nested_module (
    input logic nm_in,
    output logic nm_out
);
    assign nm_out = nm_in;
endmodule

