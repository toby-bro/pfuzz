module Module_IfNoneParam (
    input int in_port,
    output int out_port
);
    assign out_port = in_port;
endmodule

