module CoverageHelper (
    input bit in_h,
    output logic out_h
);
    assign out_h = in_h;
endmodule

